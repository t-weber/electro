../../display/sevenseg_multi.sv