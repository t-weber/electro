../lib/sevenseg.sv