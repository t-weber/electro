../../display/pixlcd_3wire.sv