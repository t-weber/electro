../../comm/serial.sv