../../clock/clkgen.sv