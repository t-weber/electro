../../display/sevenseg.sv