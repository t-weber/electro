../../display/lcd_3wire.sv