../../display/txtlcd_3wire.sv